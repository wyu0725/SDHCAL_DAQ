library verilog;
use verilog.vl_types.all;
entity DaqSwitcher is
    port(
        DaqSelect       : in     vl_logic;
        AutoDaq_PWR_ON_A: in     vl_logic;
        AutoDaq_PWR_ON_D: in     vl_logic;
        AutoDaq_PWR_ON_ADC: in     vl_logic;
        AutoDaq_PWR_ON_DAC: in     vl_logic;
        SlaveDaq_PWR_ON_A: in     vl_logic;
        SlaveDaq_PWR_ON_D: in     vl_logic;
        SlaveDaq_PWR_ON_ADC: in     vl_logic;
        SlaveDaq_PWR_ON_DAC: in     vl_logic;
        PWR_ON_D        : out    vl_logic;
        PWR_ON_A        : out    vl_logic;
        PWR_ON_ADC      : out    vl_logic;
        PWR_ON_DAC      : out    vl_logic;
        AutoDaq_RESET_B : in     vl_logic;
        SlaveDaq_RESET_B: in     vl_logic;
        RESET_B         : out    vl_logic;
        AutoDaq_START_ACQ: in     vl_logic;
        SlaveDaq_START_ACQ: in     vl_logic;
        START_ACQ       : out    vl_logic;
        CHIPSATB        : in     vl_logic;
        AutoDaq_CHIPSATB: out    vl_logic;
        SlaveDaq_CHIPSATB: out    vl_logic;
        UsbAcqStart     : in     vl_logic;
        AutoDaq_Start   : out    vl_logic;
        SlaveDaq_Start  : out    vl_logic;
        AutoDaq_StartReadout: in     vl_logic;
        SlaveDaq_StartReadout: in     vl_logic;
        StartReadout    : out    vl_logic;
        EndReadout      : in     vl_logic;
        AutoDaq_EndReadout: out    vl_logic;
        SlaveDaq_EndReadout: out    vl_logic;
        AutoDaq_OnceEnd : in     vl_logic;
        SlaveDaq_OnceEnd: in     vl_logic;
        OnceEnd         : out    vl_logic;
        AutoDaq_AllDone : in     vl_logic;
        SlaveDaq_AllDone: in     vl_logic;
        AllDone         : out    vl_logic;
        DataTransmitDone: in     vl_logic;
        AutoDaq_DataTransmitDone: out    vl_logic;
        SlaveDaq_DataTransmitDone: out    vl_logic;
        ExternalTrigger : in     vl_logic;
        SingleStart     : out    vl_logic;
        AutoDaq_UsbStartStop: in     vl_logic;
        SlaveDaq_UsbStartStop: in     vl_logic;
        UsbStartStop    : out    vl_logic
    );
end DaqSwitcher;
