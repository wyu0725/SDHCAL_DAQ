`timescale 1ns/1ns
module SCurve_Data_FIFO_tb;
reg clk;
reg rst;
reg [15:0] din;
reg wr_en;
reg rd_en;
wire [15:0] dout;
wire full;
wire empty;
SCurve_Data_FIFO uut(
  .clk(clk),
  .rst(rst),
  .din(din),
  .wr_en(wr_en),
  .rd_en(rd_en),
  .dout(dout),
  .full(full),
  .empty(empty)
);
parameter PEROID = 25;
initial begin
  clk = 1'b0;
  rst = 1'b1;
  din = 16'b0;
  wr_en = 1'b0;
  rd_en = 1'b0;
  #100;
  rst = 1'b0;
  #13;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h0;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h1;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h2;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h3;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h4;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h5;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h6;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h7;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h8;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h9;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'ha;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'hb;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'hc;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'hd;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'he;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'hf;
  #(PEROID);
  wr_en = 1'b0;
  //read
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  #(PEROID);
  rd_en = 1'b1;
  #(PEROID); 
  rd_en = 1'b0;
  //write while read
  #(PEROID);
  wr_en = 1'b1;
  din = 16'h5;
  #(PEROID);
  wr_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'ha;
  rd_en = 1'b1;
  #(PEROID);
  wr_en = 1'b0;
  rd_en = 1'b0;
  #(PEROID);
  wr_en = 1'b1;
  din = 16'hf;
  rd_en = 1'b1;
  #(PEROID);
  wr_en = 1'b0;
  rd_en = 1'b0;
end
//Generate clk
localparam High = 12;
localparam Low = 13;
always begin
  #(Low) clk = ~clk;
  #(High) clk = ~clk;
end
endmodule
