library verilog;
use verilog.vl_types.all;
entity ACQ_or_SCTest_Switch_tb is
end ACQ_or_SCTest_Switch_tb;
