`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/05/21 10:57:19
// Design Name:
// Module Name: FPGA_Top
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////
//																//
//                                                    `:/+:		//
//                                                 .odNmydMs	//
//                                               :hMNy: `dMh	//
//     ./+oo+-   -://////+oo`  `:/ooso/`       :dMNy.  .dMm-	//
//   /dNy/:/hM/ odyNMmssso+. +dNNd+/+yMM/    .hMMh- ..oNMd-		//
// `hMd-     -  ` .MMo      -m+sMN-   mMy   /NMN+ .yMMMNs`		//	
// yMm.         `ymMMmddd+  .- dMd` -hMh.  yMMd- :NMMNy.		//	
// NMh          .:NMh...`   .ymMMmdmds:   yMMm.  /dd+.    `		//
// dMm.    `+h`  :MM/         yMm-`      :MMN/         `oh-		//
// .hMNysydNd+   /MMdyyhdd`  `NMs        sMMN.       :yd+`		//
//   ./++/:.      ./++/:-`   -mm:        /MMMh:..-+ymd/`		//
//                                        +mMMMMMNdo-			//
//                                          .:/:-`				//
//																//
//////////////////////////////////////////////////////////////////
module FPGA_Top(
	input Clk40M,
	input rst_n
	);
	MicrorocControl MicrororChain1(
		);
endmodule
