library verilog;
use verilog.vl_types.all;
entity Switcher_tb is
end Switcher_tb;
