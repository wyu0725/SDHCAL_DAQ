library verilog;
use verilog.vl_types.all;
entity Switcher is
    port(
        ModeSelect      : in     vl_logic_vector(1 downto 0);
        UsbMicroroc10BitDac0: in     vl_logic_vector(9 downto 0);
        UsbMicroroc10BitDac1: in     vl_logic_vector(9 downto 0);
        UsbMicroroc10BitDac2: in     vl_logic_vector(9 downto 0);
        SCTest10BitDac  : in     vl_logic_vector(9 downto 0);
        SweepAcq10BitDac: in     vl_logic_vector(9 downto 0);
        SweepAcqDacSelect: in     vl_logic_vector(1 downto 0);
        OutMicroroc10BitDac0: out    vl_logic_vector(9 downto 0);
        OutMicroroc10BitDac1: out    vl_logic_vector(9 downto 0);
        OutMicroroc10BitDac2: out    vl_logic_vector(9 downto 0);
        UsbMicrorocChannelMask: in     vl_logic_vector(191 downto 0);
        SCTestMicrorocChannelMask: in     vl_logic_vector(191 downto 0);
        OutMicrorocChannelMask: out    vl_logic_vector(191 downto 0);
        UsbMicrorocCTestChannel: in     vl_logic_vector(63 downto 0);
        SCTestMicrorocCTestChannel: in     vl_logic_vector(63 downto 0);
        OutMicrorocCTestChannel: out    vl_logic_vector(63 downto 0);
        UsbMicrorocSCParameterLoad: in     vl_logic;
        SCTestMicrorocSCParameterLoad: in     vl_logic;
        SweepAcqMicrorocSCParameterLoad: in     vl_logic;
        OutMicrorocSCParameterLoad: out    vl_logic;
        UsbSCOrReadreg  : in     vl_logic;
        OutMicrorocSCOrReadreg: out    vl_logic;
        UsbMicrorocAcqStartStop: in     vl_logic;
        UsbSweepTestStartStop: in     vl_logic;
        OutSCTestStartStop: out    vl_logic;
        OutSweepAcqStartStop: out    vl_logic;
        SCTestDone      : in     vl_logic;
        SweepAcqDone    : in     vl_logic;
        SweepTestDone   : out    vl_logic;
        SweepTestUsbStartStop: in     vl_logic;
        OutUsbStartStop : out    vl_logic;
        SweepAcqMicrorocAcqStartStop: in     vl_logic;
        MicrorocAcqStartStop: out    vl_logic;
        MicrorocAcqData : in     vl_logic_vector(15 downto 0);
        MicrorocAcqData_en: in     vl_logic;
        SweepAcqData    : in     vl_logic_vector(15 downto 0);
        SweepAcqData_en : in     vl_logic;
        SCTestData      : in     vl_logic_vector(15 downto 0);
        SCTestData_en   : in     vl_logic;
        UsbFifoData     : out    vl_logic_vector(15 downto 0);
        UsbFifoData_en  : out    vl_logic;
        ParallelData    : out    vl_logic_vector(15 downto 0);
        ParallelData_en : out    vl_logic
    );
end Switcher;
