library verilog;
use verilog.vl_types.all;
entity SweepACQ_Control_tb is
end SweepACQ_Control_tb;
