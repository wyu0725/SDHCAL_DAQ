// Verilog created by ORCAD Capture

module PAD30X30V2 
 ( 
		GEM_OUT_A );

output	[1:64]	GEM_OUT_A;

initial
	begin
	end

endmodule
