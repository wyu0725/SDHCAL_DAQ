// Verilog created by ORCAD Capture

module PAD30X30V2 
 ( 
		GEM_OUT_I, 
		GEM_SIGNAL_S3, 
		GEM_OUT_E, 
		GEM_SIGNAL_J2, 
		GEM_OUT_L, 
		GEM_SIGNAL_S27, 
		GEM_OUT_J, 
		GEM_SIGNAL_S11, 
		GEM_OUT_O, 
		GEM_SIGNAL_AF20, 
		GEM_OUT_A, 
		GEM_SIGNAL_B4, 
		GEM_OUT_F, 
		GEM_SIGNAL_J10, 
		GEM_OUT_H, 
		GEM_SIGNAL_J26, 
		GEM_OUT_K, 
		GEM_SIGNAL_S19, 
		GEM_OUT_N, 
		GEM_SIGNAL_AF12, 
		GEM_OUT_B, 
		GEM_SIGNAL_A15, 
		GEM_OUT_D, 
		GEM_SIGNAL_D28, 
		GEM_OUT_G, 
		GEM_SIGNAL_J18, 
		GEM_OUT_M, 
		GEM_SIGNAL_AF4, 
		GEM_OUT_C, 
		GEM_SIGNAL_A23, 
		GEM_OUT_P, 
		GEM_SIGNAL_AF28 );

output	GEM_SIGNAL_S3;
output	[1:64]	GEM_OUT_I;
output	GEM_SIGNAL_J2;
output	[1:64]	GEM_OUT_E;
output	GEM_SIGNAL_S27;
output	[1:64]	GEM_OUT_L;
output	GEM_SIGNAL_S11;
output	[1:64]	GEM_OUT_J;
output	GEM_SIGNAL_AF20;
output	[1:64]	GEM_OUT_O;
output	GEM_SIGNAL_B4;
output	[1:64]	GEM_OUT_A;
output	GEM_SIGNAL_J10;
output	[1:64]	GEM_OUT_F;
output	GEM_SIGNAL_J26;
output	[1:64]	GEM_OUT_H;
output	GEM_SIGNAL_S19;
output	[1:64]	GEM_OUT_K;
output	GEM_SIGNAL_AF12;
output	[1:64]	GEM_OUT_N;
output	GEM_SIGNAL_A15;
output	[1:64]	GEM_OUT_B;
output	GEM_SIGNAL_D28;
output	[1:64]	GEM_OUT_D;
output	GEM_SIGNAL_J18;
output	[1:64]	GEM_OUT_G;
output	GEM_SIGNAL_AF4;
output	[1:64]	GEM_OUT_M;
output	GEM_SIGNAL_A23;
output	[1:64]	GEM_OUT_C;
output	GEM_SIGNAL_AF28;
output	[1:64]	GEM_OUT_P;

initial
	begin
	end

endmodule
