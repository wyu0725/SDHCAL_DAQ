// Verilog created by ORCAD Capture

module XC7A100TFGG484 
 ( 
		VMGTAVCC, 
		VMGTAVTT, 
		\SFP_RX+ , 
		GND, 
		SFP_CLK_P, 
		SFP_CLK_N, 
		\SFP_RX- , 
		\SFP_TX+ , 
		\SFP_TX- , 
		\VCC3.3VD , 
		REGULARIO_SFP_TX_DISABLE, 
		TRIGEXT_E, 
		REGULARIO_SFP_SDA, 
		CDR_SDA, 
		STARTREADOUT2_E, 
		DOUT1B_E, 
		CHIPSATB_E, 
		CDR_SCK, 
		TRANSMITON1B_E, 
		SR_CK_E, 
		SR_RSTB_E, 
		ENDREADOUT2_E, 
		REGULARIO_SFP_SCL, 
		DOUT2B_E, 
		STARTREADOUT1_E, 
		SR_IN_E, 
		STARTACQ_E, 
		TRANSMITON2B_E, 
		TRIGEXT_D, 
		TRANSMITON1B_D, 
		ENDREADOUT1_E, 
		SR_OUT_E, 
		STARTACQ_D, 
		\RESET# , 
		SR_IN_D, 
		STARTREADOUT1_D, 
		DOUT2B_D, 
		CDR_LOL, 
		SR_CK_D, 
		STARTREADOUT2_D, 
		DOUT1B_D, 
		CHIPSATB_D, 
		SR_OUT_D, 
		ENDREADOUT1_D, 
		SR_RSTB_D, 
		TRANSMITON2B_D, 
		PWR_ON_A, 
		PWR_ON_ADC, 
		PWR_ON_DAC, 
		ENDREADOUT2_D, 
		DOUT1B_C, 
		TRIGEXT_C, 
		STARTACQ_C, 
		PWR_ON_D, 
		STARTREADOUT2_C, 
		CHIPSATB_C, 
		TRANSMITON1B_C, 
		\VCC3.3VD , 
		CHIPSATB_A, 
		TRANSMITON2B_A, 
		SR_CK_A, 
		SR_OUT_A, 
		STARTREADOUT2_A, 
		OUT_TRIG1B, 
		ROWSELECT0, 
		ENDREADOUT1_A, 
		CALI_SW_A, 
		ROWSELECT1, 
		\CALI_CS# , 
		CALI_SW_B, 
		OUT_TRIG2B, 
		ADC_CLK, 
		COLUMNSELECT1, 
		ADC_DATA3, 
		ADC_DATA1, 
		ADC_DATA2, 
		ADC_DATA0, 
		TP0, 
		COLUMNSELECT2, 
		ROWSELECT2, 
		COLUMNSELECT0, 
		ENDREADOUT2_A, 
		CALI_DIN, 
		SR_IN_A, 
		SR_RSTB_A, 
		CALI_SCK, 
		DOUT2B_A, 
		STARTREADOUT1_A, 
		\VCC3.3VD , 
		DONE, 
		TCK, 
		GND, 
		VCCADC, 
		CCLK, 
		TDO, 
		TDI, 
		INIT_B, 
		TMS, 
		PROGRAM_B, 
		\VCC3.3VD , 
		SFP_TX_DISABLE, 
		FD, 
		FIFOADR0, 
		PKTEND, 
		FIFOADR1, 
		FLAGB, 
		SLOE, 
		SFP_SCL, 
		SFP_SDA, 
		FLAGA, 
		FLAGC, 
		SLWR, 
		SLRD, 
		CLKOUT, 
		CLK_40M, 
		SLCS, 
		IFCLK, 
		DTCC_DATA2OUT, 
		DTCC_CONTROL2IN, 
		DTCC_CONTROL1IN, 
		PLUG1DATAOUT1, 
		PLUG2_DATAIN1, 
		PLUG2_DATAIN2, 
		DTCC_DATA1OUT, 
		\VCC2.5VD , 
		\REGULARIO_SFP_TX+ , 
		\REGULARIO_SFP_TX- , 
		RX_CDR_RXP, 
		RX_CDR_RXN, 
		RAZ_CHNP, 
		RAZ_CHNN, 
		VAL_EVTP, 
		VAL_EVTN, 
		CK_5P, 
		CK_5N, 
		RX_CDR_CLKP, 
		RX_CDR_CLKN, 
		SPARE_LVDS_P, 
		SPARE_LVDS_N, 
		CK_40P, 
		CK_40N, 
		\VCC3.3VD , 
		TRANSMITON2B_C, 
		D00, 
		D01, 
		D02, 
		D03, 
		PUDC_B, 
		SR_CK_C, 
		SR_OUT_C, 
		STARTREADOUT1_C, 
		SR_RSTB_C, 
		FCS_B, 
		ENDREADOUT2_C, 
		ENDREADOUT1_C, 
		SELECT, 
		SR_IN_B, 
		TRANSMITON1B_B, 
		HOLD, 
		DOUT2B_B, 
		CHIPSATB_B, 
		STARTREADOUT2_B, 
		RST_COUNTERB, 
		TRIGEXT_B, 
		STARTREADOUT1_B, 
		SR_CK_B, 
		SR_OUT_B, 
		STARTACQ_A, 
		STARTACQ_B, 
		DOUT1B_B, 
		TRIGEXT_A, 
		ENDREADOUT2_B, 
		ENDREADOUT1_B, 
		TRANSMITON2B_B, 
		DOUT1B_A, 
		TRANSMITON1B_A, 
		SR_RSTB_B, 
		RESET_B, 
		OUT_TRIG0B, 
		SR_IN_C, 
		DOUT2B_C, 
		\VCC3.3VD , 
		DTCC_CLK2OUT, 
		DTCC_CLK1OUT, 
		PLUG2_CC1, 
		PLUG2_CC2, 
		PLUG1DATAOUT2, 
		PLUG1_CC2, 
		ELINKDATAOUT, 
		PLUG1_CC1, 
		ELINKDATAIN, 
		EXT_TRIG_IN, 
		LED, 
		OTR, 
		ADC_DATA, 
		ELINKCLKIN, 
		EXT_CLK_IN, 
		DTCC_CLK2IN, 
		DTCC_CLK1IN, 
		TP, 
		EXT_TRIG_OUT );

inout	VMGTAVCC, VMGTAVTT, \SFP_RX+ , GND, SFP_CLK_P, SFP_CLK_N, \SFP_RX- , \SFP_TX+ , \SFP_TX- ;
inout	\VCC3.3VD , REGULARIO_SFP_TX_DISABLE, TRIGEXT_E, REGULARIO_SFP_SDA, CDR_SDA, STARTREADOUT2_E, DOUT1B_E, CHIPSATB_E, CDR_SCK, TRANSMITON1B_E, SR_CK_E, SR_RSTB_E, ENDREADOUT2_E, REGULARIO_SFP_SCL, DOUT2B_E, STARTREADOUT1_E, SR_IN_E, STARTACQ_E, TRANSMITON2B_E, TRIGEXT_D, TRANSMITON1B_D, ENDREADOUT1_E, SR_OUT_E, STARTACQ_D, \RESET# , SR_IN_D, STARTREADOUT1_D, DOUT2B_D, CDR_LOL, SR_CK_D, STARTREADOUT2_D, DOUT1B_D, CHIPSATB_D, SR_OUT_D, ENDREADOUT1_D, SR_RSTB_D, TRANSMITON2B_D, PWR_ON_A, PWR_ON_ADC, PWR_ON_DAC, ENDREADOUT2_D, DOUT1B_C, TRIGEXT_C, STARTACQ_C, PWR_ON_D, STARTREADOUT2_C, CHIPSATB_C, TRANSMITON1B_C;
inout	\VCC3.3VD , CHIPSATB_A, TRANSMITON2B_A, SR_CK_A, SR_OUT_A, STARTREADOUT2_A, OUT_TRIG1B, ROWSELECT0, ENDREADOUT1_A, CALI_SW_A, ROWSELECT1, \CALI_CS# , CALI_SW_B, OUT_TRIG2B, ADC_CLK, COLUMNSELECT1, ADC_DATA3, ADC_DATA1, ADC_DATA2, ADC_DATA0, TP0, COLUMNSELECT2, ROWSELECT2, COLUMNSELECT0, ENDREADOUT2_A, CALI_DIN, SR_IN_A, SR_RSTB_A, CALI_SCK, DOUT2B_A, STARTREADOUT1_A;
inout	\VCC3.3VD , DONE, TCK, GND, VCCADC, CCLK, TDO, TDI, INIT_B, TMS, PROGRAM_B;
inout	\VCC3.3VD , SFP_TX_DISABLE, FIFOADR0, PKTEND, FIFOADR1, FLAGB, SLOE, SFP_SCL, SFP_SDA, FLAGA, FLAGC, SLWR, SLRD, CLKOUT, CLK_40M, SLCS, IFCLK, DTCC_DATA2OUT, DTCC_CONTROL2IN, DTCC_CONTROL1IN, PLUG1DATAOUT1, PLUG2_DATAIN1, PLUG2_DATAIN2, DTCC_DATA1OUT;
inout	[15:0]	FD;
inout	\VCC2.5VD , \REGULARIO_SFP_TX+ , \REGULARIO_SFP_TX- , RX_CDR_RXP, RX_CDR_RXN, RAZ_CHNP, RAZ_CHNN, VAL_EVTP, VAL_EVTN, CK_5P, CK_5N, RX_CDR_CLKP, RX_CDR_CLKN, SPARE_LVDS_P, SPARE_LVDS_N, CK_40P, CK_40N;
inout	\VCC3.3VD , TRANSMITON2B_C, D00, D01, D02, D03, PUDC_B, SR_CK_C, SR_OUT_C, STARTREADOUT1_C, SR_RSTB_C, FCS_B, ENDREADOUT2_C, ENDREADOUT1_C, SELECT, SR_IN_B, TRANSMITON1B_B, HOLD, DOUT2B_B, CHIPSATB_B, STARTREADOUT2_B, RST_COUNTERB, TRIGEXT_B, STARTREADOUT1_B, SR_CK_B, SR_OUT_B, STARTACQ_A, STARTACQ_B, DOUT1B_B, TRIGEXT_A, ENDREADOUT2_B, ENDREADOUT1_B, TRANSMITON2B_B, DOUT1B_A, TRANSMITON1B_A, SR_RSTB_B, RESET_B, OUT_TRIG0B, SR_IN_C, DOUT2B_C;
inout	\VCC3.3VD , DTCC_CLK2OUT, DTCC_CLK1OUT, PLUG2_CC1, PLUG2_CC2, PLUG1DATAOUT2, PLUG1_CC2, ELINKDATAOUT, PLUG1_CC1, ELINKDATAIN, EXT_TRIG_IN, OTR, ELINKCLKIN, EXT_CLK_IN, DTCC_CLK2IN, DTCC_CLK1IN, EXT_TRIG_OUT;
inout	[7:0]	LED;
inout	[11:0]	ADC_DATA;
inout	[3:0]	TP;

initial
	begin
	end

endmodule
