library verilog;
use verilog.vl_types.all;
entity DaqControl_tb is
end DaqControl_tb;
