library verilog;
use verilog.vl_types.all;
entity SCurve_Test_Top_tb is
end SCurve_Test_Top_tb;
