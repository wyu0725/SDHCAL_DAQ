library verilog;
use verilog.vl_types.all;
entity SCurve_Test_Control_tb is
end SCurve_Test_Control_tb;
