library verilog;
use verilog.vl_types.all;
entity ADC_AD9220_tb is
end ADC_AD9220_tb;
