library verilog;
use verilog.vl_types.all;
entity AdcControl_tb is
end AdcControl_tb;
