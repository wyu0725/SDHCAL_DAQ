library verilog;
use verilog.vl_types.all;
entity SweepACQ_Top_tb is
end SweepACQ_Top_tb;
